module practice_1(C,HEX0);

input [3:0]C;
output [6:0]HEX0;

assign HEX0[0] = 1;
assign HEX0[1] = 1;
assign HEX0[2] = 1;
assign HEX0[3] = 1;
assign HEX0[4] = 1;
assign HEX0[5] = 1;
assign HEX0[6] = 1;

endmodule